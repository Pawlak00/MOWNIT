R 0 1 1
R 0 3 1
V 4 0 1
R 2 3 1
R 1 3 1
R 4 2 1